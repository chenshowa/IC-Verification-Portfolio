//Packages

`include "apb_mem.sv"
`include "ahb_trans.sv"
`include "ahb_seq.sv"
`include "ahb_seqr.sv"
`include "ahb_drv.sv"
`include "ahb_monitor.sv"
`include "ahb_agent.sv"
`include "apb_trans.sv"
`include "apb_seq.sv"
`include "apb_seqr.sv"
`include "apb_drv.sv"
`include "apb_monitor.sv"
`include "apb_agent.sv"
`include "coverage.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "assertion.sv"