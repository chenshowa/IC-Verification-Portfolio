//definitions 

`define burst_size 6

`define ADDR_WIDTH  32
`define DATA_WIDTH  32